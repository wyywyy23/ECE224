* FILE: no_name.sp

********************** begin header *****************************

* Sample Spice Header file for Generic 2.5V 0.25 um process (mmi25)

.OPTIONS post NOMOD post_version=9601

**################################################
* Only Typical/Typical spice models included
.include '${MMI_TOOLS}/sue/schematics/mspice/mmi25.mod'
* NOTE: these are contrived spice models
**################################################

.param  arean(w,sdd) = '(w*sdd*1p)'
.param  areap(w,sdd) = '(w*sdd*1p)'
* Setup either one or the other of the following
* For ACM=0,2,10,12 fet models
.param  perin(w,sdd) = '(2u*(w+sdd))'
.param  perip(w,sdd) = '(2u*(w+sdd))'
* For ACM=3,13 fet models
*.param  perin(w,sdd) = '(1u*(w+2*sdd))'
*.param  perip(w,sdd) = '(1u*(w+2*sdd))'

.param ln_min   =  0.24u
.param lp_min   =  0.24u

* used in source/drain area/perimeter calculation
.param sdd        =  0.66

.PARAM vddp=2.25	$ VDD voltage

VDD vdd 0 DC vddp 

.TEMP 105
.TRAN 5p 10n

*********************** end header ******************************

* SPICE netlist for "no_name" generated by MMI_SUE5.6.11 on Sat Apr 16 
*+ 16:02:32 PDT 2016.

* start main CELL no_name
* .SUBCKT no_name  
X_1 out in gnd gnd enm W=1 L=ln_min ad='arean(1,sdd)' as='arean(1,sdd)' 
+ pd='perin(1,sdd)' ps='perin(1,sdd)' 
X_2 out in vdd vdd epm W='2' L=lp_min ad='areap(2,sdd)' 
+ as='areap(2,sdd)' pd='perip(2,sdd)' ps='perip(2,sdd)' 
Vvin in gnd DC 5V 
* .ENDS	$ no_name

.GLOBAL gnd vdd

.END

